module mp4datapath
(

);



endmodule mp4datapath