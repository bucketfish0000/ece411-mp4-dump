module dec_exe_reg(

)

endmodule:dec_exe_reg