module stage_fetch
(
    
);

endmodule stage_fetch