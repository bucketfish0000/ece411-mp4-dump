module fet_dec_reg
    import rv32i_types::*;
    import immediates::*; 
(
    input logic clk,
    input logic rst,
    input logic if_de_rst,
    input logic load,
    input logic sp_ld_commit,
    input logic ld_commit,

    input logic ready_i,
    output logic ready_o,
    output logic valid_o,

    input rv32i_word instr_fetch,
    input rv32i_word pc_fetch,
    input rv32i_word pc_wdata,

    output rv32i_word instr_decode,
    output rv32i_word pc_decode,
    output rv32i_word pc_wdata_decode,

    output logic [63:0] commit_order
);

    logic ready;
    logic[31:0] instr,pc_r, pc_w;
    logic [63:0] order_counter;

    always_ff @(posedge clk)
    begin
        if (rst || if_de_rst)
        begin
            ready<='0;
            instr<=0;
            pc_r<=0;
            pc_w<=0;
        end
        else if (load)
        begin
            ready<=ready_i;
            instr<=instr_fetch;
            pc_r<=pc_fetch;
            pc_w<=pc_wdata;
        end
    end
    
    always_ff @( posedge clk, posedge rst ) begin : counter_reg
        if(rst)
            order_counter <= 64'hffffffffffffffff;
        else if((load||ld_commit) && !if_de_rst)
            order_counter <= order_counter + 64'b01;
        else if(if_de_rst && sp_ld_commit) begin
            //min 4800 clk cycle, 1.28e+04 power draw, shaves 5.5 seconds off of 10000 cycle time
            order_counter <= order_counter - 64'b01;
            //if we cheat we can get to clock cycle of 4400, maybe a bit lower. Assumes that only bottom 24 bits will be used
            //saves like 5.5 seconds in coremark im vs 4800 clk cycle, but 1.38e+04 power draw
            // order_counter <= {40'h0, order_counter[23:0] - 24'b01};
        end
    end

    always_comb
    begin
        ready_o=ready;
        instr_decode=instr;
        pc_decode=pc_r;
        pc_wdata_decode=pc_w;
        commit_order = order_counter; 
    end

    //valid register
    always_ff @(posedge clk, posedge rst) begin : valid_reg
        if(rst) begin
            valid_o <= 1'b0;
        end
        else if(if_de_rst) begin
            valid_o <= 1'b0;
        end
        else if((load == 1)) begin
            valid_o <= 1'b1;
        end
    end
endmodule : fet_dec_reg

module dec_exe_reg
    import rv32i_types::*;
    import hazards::*;
    import cpuIO::*;
(
    input logic clk,
    input logic rst,
    input logic load,
    input immediates::imm imm_in,

    output immediates::imm imm_out,

    input logic ready_i,
    output logic ready_o,
    output logic valid_o,
    input rv32i_opcode opcode_dec,
    output rv32i_opcode opcode_dec_exe,

    input control_word cw_in,
    output control_word cw_out,

    output hzds instruct_in_exe
);

    immediates::imm imm_data;
    logic ready;
    control_word cw_data;
    rv32i_opcode opcode_data;
    always_ff @(posedge clk)
    begin
        if (rst) begin

            imm_data.i_imm <= 32'b0;
            imm_data.u_imm <= 32'b0;
            imm_data.b_imm <= 32'b0;
            imm_data.s_imm <= 32'b0;
            imm_data.j_imm <= 32'b0;
            opcode_data<= rv32i_opcode'(7'b0);
            ready<= 1'b0;

            cw_data.exe.cmp_sel <= cmpmux::rs2_out;
            cw_data.exe.alumux1_sel <= alumux::rs1_out;
            cw_data.exe.alumux2_sel <= alumux::i_imm;
            cw_data.exe.rs1_sel <= rs1mux::rs1_data;
            cw_data.exe.rs2_sel <= rs2mux::rs2_data;
            cw_data.exe.cmpop <= beq;
            cw_data.exe.aluop <= alu_add;
            cw_data.exe.exefwdmux_sel <= exefwdmux::alu_out;
            cw_data.exe.rs1signunsignmux_sel <= rs1signunsignmux::sign;
            cw_data.exe.rs2signunsignmux_sel <= rs2signunsignmux::sign;
            cw_data.exe.multihighlowmux_sel <= multihighlowmux::low;
            cw_data.exe.divremquotmux_sel <= divremquotmux::quotient;
            cw_data.mem.mem_read_d <= 1'b0;
            cw_data.mem.mem_write_d <= 1'b0;
            cw_data.mem.store_funct3 <= sb;
            cw_data.mem.load_funct3 <= lb;
            cw_data.mem.mar_sel <= marmux::pc_out;
            cw_data.mem.memfwdmux_sel <= memfwdmux::mem_fwd_data;
            cw_data.wb.ld_reg <= 1'b0;
            cw_data.wb.regfilemux_sel <= regfilemux::alu_out;
            cw_data.wb.rd_sel <= 5'b00000;
            cw_data.rvfi.valid_commit <= 1'b0;//done
            cw_data.rvfi.order_commit <= 64'b0;//done
            cw_data.rvfi.instruction <= 32'b0;//done
            cw_data.rvfi.rs1_addr <= 5'b0; //done
            cw_data.rvfi.rs2_addr <= 5'b0; //dome
            cw_data.rvfi.rs1_data <= 32'b0; //done
            cw_data.rvfi.rs2_data <= 32'b0; //done
            cw_data.rvfi.rd_wdata <= 32'b0;//done
            cw_data.rvfi.pc_rdata <= 32'h40000000;//done
            cw_data.rvfi.pc_wdata <= 32'b0;//done
            cw_data.rvfi.mem_addr <= 32'b0;//done
            cw_data.rvfi.rmask <= 4'b0;//done
            cw_data.rvfi.wmask <= 4'b0;//done
            cw_data.rvfi.mem_rdata <= 32'b0;//done
            cw_data.rvfi.mem_wdata <= 32'b0;//done
        end
        else if (load) begin
            imm_data<=imm_in;
            ready<=ready_i;
            opcode_data <= opcode_dec;
            cw_data<=cw_in;
        end
    end 

    always_comb
    begin
        imm_out=imm_data;
        ready_o = ready;
        cw_out=cw_data;
        opcode_dec_exe=rv32i_opcode'(cw_data.rvfi.instruction[6:0]);
    end

    always_comb begin : hzd_reg_in_exe
        instruct_in_exe.opcode = rv32i_opcode'(cw_data.rvfi.instruction[6:0]);
        instruct_in_exe.rd_addr = cw_data.wb.rd_sel;
        instruct_in_exe.rs1_addr = cw_data.rvfi.rs1_addr;
        instruct_in_exe.rs2_addr = cw_data.rvfi.rs2_addr;
        instruct_in_exe.commit_order = cw_data.rvfi.order_commit;
    end

    //valid register
    always_ff @(posedge clk) begin : valid_reg
        if(rst) begin
            valid_o <= 1'b0;
        end
        else if((load == 1)) begin
            valid_o <= 1'b1;
        end
    end

endmodule : dec_exe_reg

//substantially more complicated than other registers on account of needing to prime mar/mdo/mem_data_out for mem_stage to then be able to 
//start r/w right away
module exe_mem_reg
// Mux types are in their own packages to prevent identiier collisions
// e.g. pcmux::pc_plus4 and regfilemux::pc_plus4 are seperate identifiers
// for seperate enumerated types, you cannot //import rv32i_mux_types::*;
import rv32i_types::*;
import hazards::*;
import cpuIO::*;
(
    input logic clk, //from datapath
    input logic rst, //from datapath
    input logic exe_mem_rst,

    input logic br_en_i, 
    input logic exe_mem_ld, 
    input logic exe_rdy,
    input logic [31:0] alu_out_i,
    input logic [31:0] rs1_out_i, 
    input logic [31:0] rs2_out_i,
    input logic [31:0] u_imm_i, 

    output logic [31:0] exe_fwd_data, 
    output logic [31:0] u_imm_o, 
    output logic br_en_o, 
    output logic exe_mem_valid, 
    output logic exe_mem_rdy, 

    output logic [31:0] mem_address_d, //to data cache
    output logic [31:0] mem_wdata_d, //to data cache
    output logic [3:0] mem_byte_enable, //to data cache

    input control_word cw_in,
    output control_word cw_out,

    output logic [3:0] wmask,

    output hzds instruct_in_mem
);

    logic [31:0] fwd_temp;
    control_word cw_data;
    logic[31:0] rs2_to_mem;

    logic [31:0] marmux_o, mem_addr;
    logic trap;
    logic [3:0] rmask, wmask_temp;

    always_comb begin : exe_fwd_mux
        unique case(cw_in.exe.exefwdmux_sel)
            exefwdmux::alu_out: fwd_temp = alu_out_i;
            exefwdmux::br_en_zext: fwd_temp = {31'b0, br_en_i};
            exefwdmux::u_imm: fwd_temp = u_imm_i;
            exefwdmux::jalr: fwd_temp = cw_in.rvfi.pc_rdata + 32'h04;
        endcase
    end

    //serves as alu_out reg/fwding exe data reg for cp2 onward
    always_ff @ (posedge clk, posedge rst) begin : fwd_EX_reg
        if(rst)begin
            exe_fwd_data <= 32'b0;
        end
        else if((exe_mem_ld == 1)) begin
            exe_fwd_data <= fwd_temp;
        end
    end

    //control word reg 
     always_ff @ (posedge clk, posedge rst) begin : cw_register
        if(rst)begin
            cw_data.exe.cmp_sel <= cmpmux::rs2_out;
            cw_data.exe.alumux1_sel <= alumux::rs1_out;
            cw_data.exe.alumux2_sel <= alumux::i_imm;
            cw_data.exe.rs1_sel <= rs1mux::rs1_data;
            cw_data.exe.rs2_sel <= rs2mux::rs2_data;
            cw_data.exe.cmpop <= beq;
            cw_data.exe.aluop <= alu_add;
            cw_data.exe.exefwdmux_sel <= exefwdmux::alu_out;
            cw_data.exe.rs1signunsignmux_sel <= rs1signunsignmux::sign;
            cw_data.exe.rs2signunsignmux_sel <= rs2signunsignmux::sign;
            cw_data.exe.multihighlowmux_sel <= multihighlowmux::low;
            cw_data.exe.divremquotmux_sel <= divremquotmux::quotient;
            cw_data.mem.mem_read_d <= 1'b0;
            cw_data.mem.mem_write_d <= 1'b0;
            cw_data.mem.store_funct3 <= sb;
            cw_data.mem.load_funct3 <= lb;
            cw_data.mem.mar_sel <= marmux::pc_out;
            cw_data.mem.memfwdmux_sel <= memfwdmux::mem_fwd_data;
            cw_data.wb.ld_reg <= 1'b0;
            cw_data.wb.regfilemux_sel <= regfilemux::alu_out;
            cw_data.wb.rd_sel <= 5'b00000;
            cw_data.rvfi.valid_commit <= 1'b0;//done
            cw_data.rvfi.order_commit <= 64'b0;//done
            cw_data.rvfi.instruction <= 32'b0;//done
            cw_data.rvfi.rs1_addr <= 5'b0; //done
            cw_data.rvfi.rs2_addr <= 5'b0; //dome
            cw_data.rvfi.rs1_data <= 32'b0; //done
            cw_data.rvfi.rs2_data <= 32'b0; //done
            cw_data.rvfi.rd_wdata <= 32'b0;//done
            cw_data.rvfi.pc_rdata <= 32'h40000000;//done
            cw_data.rvfi.pc_wdata <= 32'b0;//done
            cw_data.rvfi.mem_addr <= 32'b0;//done
            cw_data.rvfi.rmask <= 4'b0;//done
            cw_data.rvfi.wmask <= 4'b0;//done
            cw_data.rvfi.mem_rdata <= 32'b0;//done
            cw_data.rvfi.mem_wdata <= 32'b0;//done
        end
        else if((exe_mem_ld == 1)) begin
            cw_data.exe <= cw_in.exe;
            cw_data.mem <= cw_in.mem;
            cw_data.wb <= cw_in.wb;
            cw_data.rvfi.valid_commit <= cw_in.rvfi.valid_commit;//done
            cw_data.rvfi.order_commit <= cw_in.rvfi.order_commit;//done
            cw_data.rvfi.instruction <= cw_in.rvfi.instruction;//done
            cw_data.rvfi.rs1_addr <= cw_in.rvfi.rs1_addr; //done
            cw_data.rvfi.rs2_addr <= cw_in.rvfi.rs2_addr; //dome
            cw_data.rvfi.rs1_data <= rs1_out_i; //done
            cw_data.rvfi.rs2_data <= rs2_out_i; //done
            cw_data.rvfi.rd_wdata <= cw_in.rvfi.rd_wdata;//done
            cw_data.rvfi.pc_rdata <= cw_in.rvfi.pc_rdata;//done
            cw_data.rvfi.pc_wdata <= cw_in.rvfi.pc_wdata;//done
            cw_data.rvfi.mem_addr <= mem_addr;//done
            cw_data.rvfi.rmask <= rmask;//done
            cw_data.rvfi.wmask <= wmask_temp;//done
            cw_data.rvfi.mem_rdata <= cw_in.rvfi.mem_rdata;//done
            cw_data.rvfi.mem_wdata <= rs2_to_mem;//done
        end
    end

    assign cw_out = cw_data;

    always_comb begin : hzd_reg_in_mem
        instruct_in_mem.opcode = rv32i_opcode'(cw_data.rvfi.instruction[6:0]);
        instruct_in_mem.rd_addr = cw_data.wb.rd_sel;
        instruct_in_mem.rs1_addr = cw_data.rvfi.rs1_addr;
        instruct_in_mem.rs2_addr = cw_data.rvfi.rs2_addr;
        instruct_in_mem.commit_order = cw_data.rvfi.order_commit;
    end

    //br_en register
    always_ff @ (posedge clk, posedge rst) begin : br_en_register
        if(rst)begin
            br_en_o <= 1'b0;
        end
        else if((exe_mem_ld == 1)) begin
            br_en_o <= br_en_i;
        end
    end

    //valid register
    always_ff @(posedge clk, posedge rst) begin : valid_reg
        if(rst) begin
            exe_mem_valid <= 1'b0;
        end
        else if(exe_mem_rst) begin
            exe_mem_valid <= 1'b0;
        end
        else if((exe_mem_ld == 1)) begin
            exe_mem_valid <= 1'b1;
        end
    end

    //ready register
    always_ff @(posedge clk, posedge rst) begin : ready_reg
        if(rst) begin
            exe_mem_rdy <= 1'b0;
        end
        else if((exe_mem_ld == 1)) begin
            exe_mem_rdy <= exe_rdy;
        end
    end

    //u_imm register
    always_ff @ (posedge clk, posedge rst) begin : u_imm_register
        if(rst)begin
            u_imm_o <= 32'b0;
        end
        else if((exe_mem_ld == 1)) begin
            u_imm_o <= u_imm_i;
        end
    end

    //include these here bc they need to be loaded at same time as EXE_MEM
    //also have rvfi signals here, mem_byte_enable is only able to be calculated once
    //we have address(which is only available after exe computes it)
    assign wmask = wmask_temp;

    always_comb begin : mem_mux
        unique case (cw_in.mem.mar_sel)
            marmux::pc_out: marmux_o = cw_in.rvfi.pc_rdata;
            marmux::alu_out: marmux_o = alu_out_i;
        endcase
    end

    
    always_comb begin : calc_addr
        rmask = 4'b0000;
        wmask_temp = 4'b0000;
        mem_addr = marmux_o;
        rs2_to_mem = rs2_out_i;
        trap = 1'b0;

        if(cw_in.mem.mem_read_d) begin
            case (cw_in.mem.load_funct3)
                lw: begin
                    rmask = 4'b1111;
                end
                lh, lhu: begin
                    rmask = (4'b0011) << (marmux_o%4); /* Modify for MP1 Final */ //correct???
                    mem_addr = marmux_o - (marmux_o%4);
                end
                lb, lbu: begin
                    rmask = (4'b0001) << (marmux_o%4); /* Modify for MP1 Final */ //correct???
                    mem_addr = marmux_o - (marmux_o%4);
                end
                default: trap = '1;
            endcase
        end
        else if(cw_in.mem.mem_write_d) begin
            case (cw_in.mem.store_funct3)
                sw: begin
                    wmask_temp = 4'b1111;
                end
                sh: begin
                    wmask_temp = (4'b0011) << (marmux_o%4); /* Modify for MP1 Final */ //correct???
                    mem_addr = marmux_o - (marmux_o%4);
                    rs2_to_mem = rs2_out_i << (8*(marmux_o%4));
                end
                sb: begin
                    wmask_temp = (4'b0001) << (marmux_o%4); /* Modify for MP1 Final */ //correct???
                    mem_addr = marmux_o - (marmux_o%4);
                    rs2_to_mem = rs2_out_i << (8*(marmux_o%4));
                end
                default: trap = '1;
            endcase
        end
        else begin
            //if not ld or st, don't really care what outputs are so just leave as default
        end
    end

    //mem_byte_enable register
    always_ff @ (posedge clk, posedge rst) begin : mem_byte_enable_register
        if(rst)begin
            mem_byte_enable <= 4'b0000;
        end
        else if((exe_mem_ld == 1) && ((cw_in.mem.mem_read_d) || (cw_in.mem.mem_write_d))) begin
            if(cw_in.mem.mem_read_d) begin
                mem_byte_enable <= rmask;
            end
            else if(cw_in.mem.mem_write_d) begin
                mem_byte_enable <= wmask_temp;
            end
        end
    end

    mem_data_out mdo_reg(
        .clk(clk),
        .reset(rst),
        .load_data_out((exe_mem_ld == 1) && ((cw_in.mem.mem_read_d) || (cw_in.mem.mem_write_d))),
        .mdo_in(rs2_to_mem),//fill in the shifted data: 
        .mdo_out(mem_wdata_d)
    );
    
    mar mar_reg(
        .clk(clk),
        .reset(rst),
        .load_mar((exe_mem_ld == 1) && ((cw_in.mem.mem_read_d) || (cw_in.mem.mem_write_d))),
        .mar_in(mem_addr),
        .mar_out(mem_address_d)
    );

endmodule : exe_mem_reg



module mem_wb_reg
    import rv32i_types::*;
    import hazards::*;
    import cpuIO::*;
(
    input clk,
    input rst,
    input logic mem_wb_ld,
    input logic mem_rdy,
    input logic [31:0] alu_out_i, //aka exe_fwd_data
    input logic br_en_i,
    input logic [31:0] u_imm_i,
    input logic [31:0] mem_rdata_D_i,
    output logic [31:0] u_imm_o,
    output logic [31:0] mem_rdata_D_o,
    output logic [31:0] mem_fwd_data,
    output logic mem_wb_rdy,
    output logic mem_wb_valid,
    output logic [31:0] alu_out_o, //aka exe_fwd_data
    output logic br_en_o,

    input control_word cw_in,
    output control_word cw_out,

    output hzds instruct_in_wb
);
    logic [31:0] alu_out_r, u_imm_r, mem_rdata_r, memfwdmux_o, mem_fwd_data_r, whole_byte, whole_half, true_mem_i;
    control_word cw_data;
    logic br_en_r, valid_r, ready_r;
    logic [7:0] byte_in;
    logic [15:0] half_in;

    always_comb begin : mem_data_slice_selection
        case(cw_in.rvfi.rmask)
            4'b0001: begin
                byte_in = mem_rdata_D_i[7:0];
                half_in = 16'hb00b;
            end
            4'b0010: begin
                byte_in = mem_rdata_D_i[15:8];
                half_in = 16'hb00b;
            end
            4'b0100: begin
                byte_in = mem_rdata_D_i[23:16];
                half_in = 16'hb00b;
            end
            4'b1000: begin
                byte_in = mem_rdata_D_i[31:24];
                half_in = 16'hb00b;
            end
            4'b0011: begin
                byte_in = 8'hab;
                half_in = mem_rdata_D_i[15:0];
            end
            4'b1100: begin
                byte_in = 8'hab;
                half_in = mem_rdata_D_i[31:16];
            end
            default: begin
                byte_in = 8'hab;
                half_in = 16'hb00b;
            end
        endcase
    end

    sext_byte sexy_byte(
        .byte_in(byte_in),
        .whole_byte_out(whole_byte)
    );

    sext_half sexy_half(
        .half_in(half_in),
        .whole_half_out(whole_half)
    );

    always_comb begin
        case(cw_in.wb.regfilemux_sel)
            regfilemux::lb: true_mem_i = whole_byte;
            regfilemux::lbu: true_mem_i = {24'b0, byte_in};
            regfilemux::lh: true_mem_i = whole_half;
            regfilemux::lhu: true_mem_i = {16'b0, half_in};
            default: true_mem_i = mem_rdata_D_i;
        endcase
    end

    always_comb begin : memfwdmux
        unique case(cw_in.mem.memfwdmux_sel)
            memfwdmux::mem_fwd_data: memfwdmux_o = true_mem_i;
            memfwdmux::exe_fwd_data: memfwdmux_o = alu_out_i;
            memfwdmux::pc_plus_4: memfwdmux_o = cw_in.rvfi.pc_rdata + 4;
        endcase
    end

    //mem_fwd_data reg
    always_ff @ (posedge clk, posedge rst) begin : mem_fwd_data_reg
        if(rst)begin
            mem_fwd_data <= 32'b0;
        end
        else if((mem_wb_ld == 1)) begin
            mem_fwd_data <= memfwdmux_o;
        end
    end

    //mem_rdata reg
    always_ff @ (posedge clk, posedge rst) begin : mem_rdata_reg
        if(rst)begin
            mem_rdata_D_o <= 32'b0;
        end
        else if((mem_wb_ld == 1)) begin
            mem_rdata_D_o <= true_mem_i;
        end
    end

    //serves as alu_out reg/fwding exe data reg for cp2 onward
    always_ff @ (posedge clk, posedge rst) begin : alu_out_reg
        if(rst)begin
            alu_out_o <= 32'b0;
        end
        else if((mem_wb_ld == 1)) begin
            alu_out_o <= alu_out_i;
        end
    end


    //control word for WB 
    always_ff @ (posedge clk, posedge rst) begin : cw_register
        if(rst)begin
            cw_data.exe.cmp_sel <= cmpmux::rs2_out;
            cw_data.exe.alumux1_sel <= alumux::rs1_out;
            cw_data.exe.alumux2_sel <= alumux::i_imm;
            cw_data.exe.rs1_sel <= rs1mux::rs1_data;
            cw_data.exe.rs2_sel <= rs2mux::rs2_data;
            cw_data.exe.cmpop <= beq;
            cw_data.exe.aluop <= alu_add;
            cw_data.exe.exefwdmux_sel <= exefwdmux::alu_out;
            cw_data.exe.rs1signunsignmux_sel <= rs1signunsignmux::sign;
            cw_data.exe.rs2signunsignmux_sel <= rs2signunsignmux::sign;
            cw_data.exe.multihighlowmux_sel <= multihighlowmux::low;
            cw_data.exe.divremquotmux_sel <= divremquotmux::quotient;
            cw_data.mem.mem_read_d <= 1'b0;
            cw_data.mem.mem_write_d <= 1'b0;
            cw_data.mem.store_funct3 <= sb;
            cw_data.mem.load_funct3 <= lb;
            cw_data.mem.mar_sel <= marmux::pc_out;
            cw_data.mem.memfwdmux_sel <= memfwdmux::mem_fwd_data;
            cw_data.wb.ld_reg <= 1'b0;
            cw_data.wb.regfilemux_sel <= regfilemux::alu_out;
            cw_data.wb.rd_sel <= 5'b00000;
            cw_data.rvfi.valid_commit <= 1'b0;//done
            cw_data.rvfi.order_commit <= 64'b0;//done
            cw_data.rvfi.instruction <= 32'b0;//done
            cw_data.rvfi.rs1_addr <= 5'b0; //done
            cw_data.rvfi.rs2_addr <= 5'b0; //dome
            cw_data.rvfi.rs1_data <= 32'b0; //done
            cw_data.rvfi.rs2_data <= 32'b0; //done
            cw_data.rvfi.rd_wdata <= 32'b0;//done
            cw_data.rvfi.pc_rdata <= 32'h40000000;//done
            cw_data.rvfi.pc_wdata <= 32'b0;//done
            cw_data.rvfi.mem_addr <= 32'b0;//done
            cw_data.rvfi.rmask <= 4'b0;//done
            cw_data.rvfi.wmask <= 4'b0;//done
            cw_data.rvfi.mem_rdata <= 32'b0;//done
            cw_data.rvfi.mem_wdata <= 32'b0;//done
        end
        else if((mem_wb_ld == 1)) begin
            if(cw_data.rvfi.instruction[6:0] == 7'b0000011) begin
                cw_data.exe <= cw_in.exe;
                cw_data.mem <= cw_in.mem;
                cw_data.wb <= cw_in.wb;
                cw_data.rvfi.valid_commit <= cw_in.rvfi.valid_commit;//done
                cw_data.rvfi.order_commit <= cw_in.rvfi.order_commit;//done
                cw_data.rvfi.instruction <= cw_in.rvfi.instruction;//done
                cw_data.rvfi.rs1_addr <= cw_in.rvfi.rs1_addr; //done
                cw_data.rvfi.rs2_addr <= cw_in.rvfi.rs2_addr; //dome
                cw_data.rvfi.rs1_data <= cw_in.rvfi.rs1_data; //done
                cw_data.rvfi.rs2_data <= cw_in.rvfi.rs2_data; //done
                cw_data.rvfi.rd_wdata <= true_mem_i;//done
                cw_data.rvfi.pc_rdata <= cw_in.rvfi.pc_rdata;//done
                cw_data.rvfi.pc_wdata <= cw_in.rvfi.pc_wdata;//done
                cw_data.rvfi.mem_addr <= cw_in.rvfi.mem_addr;//done
                cw_data.rvfi.rmask <= cw_in.rvfi.rmask;//done
                cw_data.rvfi.wmask <= cw_in.rvfi.wmask;//done
                cw_data.rvfi.mem_rdata <= mem_rdata_D_i;//done
                cw_data.rvfi.mem_wdata <= cw_in.rvfi.mem_wdata;//done
            end
            else begin
                cw_data.exe <= cw_in.exe;
                cw_data.mem <= cw_in.mem;
                cw_data.wb <= cw_in.wb;
                cw_data.rvfi.valid_commit <= cw_in.rvfi.valid_commit;//done
                cw_data.rvfi.order_commit <= cw_in.rvfi.order_commit;//done
                cw_data.rvfi.instruction <= cw_in.rvfi.instruction;//done
                cw_data.rvfi.rs1_addr <= cw_in.rvfi.rs1_addr; //done
                cw_data.rvfi.rs2_addr <= cw_in.rvfi.rs2_addr; //dome
                cw_data.rvfi.rs1_data <= cw_in.rvfi.rs1_data; //done
                cw_data.rvfi.rs2_data <= cw_in.rvfi.rs2_data; //done
                cw_data.rvfi.rd_wdata <= cw_in.rvfi.rd_wdata;//done
                cw_data.rvfi.pc_rdata <= cw_in.rvfi.pc_rdata;//done
                cw_data.rvfi.pc_wdata <= cw_in.rvfi.pc_wdata;//done
                cw_data.rvfi.mem_addr <= cw_in.rvfi.mem_addr;//done
                cw_data.rvfi.rmask <= cw_in.rvfi.rmask;//done
                cw_data.rvfi.wmask <= cw_in.rvfi.wmask;//done
                cw_data.rvfi.mem_rdata <= mem_rdata_D_i;//done
                cw_data.rvfi.mem_wdata <= cw_in.rvfi.mem_wdata;//done
            end
        end
    end

    assign cw_out = cw_data;

    always_comb begin : hzd_reg_in_wb
        instruct_in_wb.opcode = rv32i_opcode'(cw_data.rvfi.instruction[6:0]);
        instruct_in_wb.rd_addr = cw_data.wb.rd_sel;
        instruct_in_wb.rs1_addr = cw_data.rvfi.rs1_addr;
        instruct_in_wb.rs2_addr = cw_data.rvfi.rs2_addr;
        instruct_in_wb.commit_order = cw_data.rvfi.order_commit;
    end

    //br_en register
    always_ff @ (posedge clk, posedge rst) begin : br_en_register
        if(rst)begin
            br_en_o <= 1'b0;
        end
        else if((mem_wb_ld == 1)) begin
            br_en_o <= br_en_i;
        end
    end

    //valid register
    always_ff @(posedge clk, posedge rst) begin : valid_reg
        if(rst) begin
            mem_wb_valid <= 1'b0;
        end
        else if((mem_wb_ld == 1)) begin
            mem_wb_valid <= 1'b1;
        end
    end

    //ready register
    always_ff @(posedge clk, posedge rst) begin : ready_reg
        if(rst) begin
            mem_wb_rdy <= 1'b0;
        end
        else if((mem_wb_ld == 1)) begin
            mem_wb_rdy <= mem_rdy;
        end
    end

    //u_imm register
    always_ff @ (posedge clk, posedge rst) begin : u_imm_register
        if(rst)begin
            u_imm_o <= 32'b0;
        end
        else if((mem_wb_ld == 1)) begin
            u_imm_o <= u_imm_i;
        end
    end



endmodule : mem_wb_reg


module wb_fwd_reg(
    input clk,
    input rst,
    input load_wb_fwd_reg,
    input logic [31:0] wb_fwd_data_i,

    output logic [31:0] wb_fwd_data_o
);
    always_ff @ (posedge clk, posedge rst) begin : wb_fwd_register
        if(rst) begin
            wb_fwd_data_o <= 32'b0;
        end
        else if(load_wb_fwd_reg) begin
            wb_fwd_data_o <= wb_fwd_data_i;
        end
    end

endmodule : wb_fwd_reg
