
module control
import rv32i_types::*; /* Import types defined in rv32i_types.sv */
(
    input clk,
    input rst,
    input rv32i_opcode opcode,
    input logic [2:0] funct3,
    input logic [6:0] funct7,
    input logic br_en,
    input logic [4:0] rs1,
    input logic [4:0] rs2,
    input mem_resp, //added
    input rv32i_word mem_address, //added
    output pcmux::pcmux_sel_t pcmux_sel,
    output alumux::alumux1_sel_t alumux1_sel,
    output alumux::alumux2_sel_t alumux2_sel,
    output regfilemux::regfilemux_sel_t regfilemux_sel,
    output marmux::marmux_sel_t marmux_sel,
    output cmpmux::cmpmux_sel_t cmpmux_sel,
    output alu_ops aluop,
    output bit [2:0] cmpop, //added
    output logic load_pc,
    output logic load_ir,
    output logic load_regfile,
    output logic load_mar,
    output logic load_mdr,
    output logic load_data_out,
    output logic mem_read, //added
    output logic mem_write, //added
    output logic [3:0] mem_byte_enable, //added
    output rv32i_word mem_addr //added
);

/***************** USED BY RVFIMON --- ONLY MODIFY WHEN TOLD *****************/
logic trap;
logic [4:0] rs1_addr, rs2_addr;
logic [3:0] rmask, wmask;
/*****************************************************************************/

branch_funct3_t branch_funct3;
store_funct3_t store_funct3;
load_funct3_t load_funct3;
arith_funct3_t arith_funct3;

assign arith_funct3 = arith_funct3_t'(funct3);
assign branch_funct3 = branch_funct3_t'(funct3);
assign load_funct3 = load_funct3_t'(funct3);
assign store_funct3 = store_funct3_t'(funct3);
assign rs1_addr = rs1;
assign rs2_addr = rs2;

always_comb
begin : trap_check
    trap = '0;
    rmask = '0;
    wmask = '0;
    mem_addr = mem_address;

    case (opcode)
        op_lui: begin
            
        end
        
        op_auipc: begin
            
        end
        
        op_imm: begin
            
        end
        
        op_reg: begin
            
        end
        
        op_jal: begin
            
        end
         
        op_jalr: begin
            
        end

        op_br: begin
            case (branch_funct3)
                beq: begin
                    
                end
                bne: begin
                    
                end
                blt: begin
                    
                end
                bge: begin
                    
                end
                bltu: begin
                    
                end
                bgeu: begin
                        
                end
                default: trap = '1;
            endcase
        end

        op_load: begin
            case (load_funct3)
                lw: rmask = 4'b1111;
                lh, lhu: begin
                    rmask = (4'b0011) << (mem_address%4); /* Modify for MP1 Final */ //correct???
                    mem_addr = mem_address - (mem_address%4);
                end
                lb, lbu: begin
                    rmask = (4'b0001) << (mem_address%4); /* Modify for MP1 Final */ //correct???
                    mem_addr = mem_address - (mem_address%4);
                end
                default: trap = '1;
            endcase
        end

        op_store: begin
            case (store_funct3)
                sw: wmask = 4'b1111;
                sh: begin
                    wmask = (4'b0011) << (mem_address%4); /* Modify for MP1 Final */ //correct???
                    mem_addr = mem_address - (mem_address%4);
                end
                sb: begin
                    wmask = (4'b0001) << (mem_address%4); /* Modify for MP1 Final */ //correct???
                    mem_addr = mem_address - (mem_address%4);
                end
                default: trap = '1;
            endcase
        end

        default: trap = '1;
    endcase
end
/*****************************************************************************/

enum int unsigned { /* List of states */
    f1 = 0,
    f2 = 1,
    f3 = 2,
    de = 3,
    imm = 4,
    lui = 5,
    br = 6,
    auipc = 7,
    calc_addr = 8,
    ld1 = 9,
    ld2 = 10,
    st1 = 11,
    st2 = 12,
    reg0 = 13,
    jal = 14,
    jalr = 15
} state, next_states;

/************************* Function Definitions *******************************/
/**
 *  You do not need to use these functions, but it can be nice to encapsulate
 *  behavior in such a way.  For example, if you use the `loadRegfile`
 *  function, then you only need to ensure that you set the load_regfile bit
 *  to 1'b1 in one place, rather than in many.
 *
 *  SystemVerilog functions must take zero "simulation time" (as opposed to 
 *  tasks).  Thus, they are generally synthesizable, and appropraite
 *  for design code.  Arguments to functions are, by default, input.  But
 *  may be passed as outputs, inouts, or by reference using the `ref` keyword.
**/

/**
 *  Rather than filling up an always_block with a whole bunch of default values,
 *  set the default values for controller output signals in this function,
 *   and then call it at the beginning of your always_comb block.
**/
alu_ops alu_oppy;

function void set_defaults();
    pcmux_sel = pcmux::pc_plus4;
    alumux1_sel = alumux::rs1_out;
    alumux2_sel = alumux::i_imm;
    regfilemux_sel = regfilemux::alu_out;
    marmux_sel = marmux::pc_out;
    cmpmux_sel = cmpmux::rs2_out;
    $cast(alu_oppy, 3'b000);
    aluop = alu_oppy;
    cmpop = 3'b000;
    load_pc = 1'b0;
    load_ir = 1'b0;
    load_regfile = 1'b0;
    load_mar = 1'b0;
    load_mdr = 1'b0;
    load_data_out = 1'b0;
    mem_read = 1'b0;
    mem_write = 1'b0;
    mem_byte_enable = 4'b1111;
endfunction

/**
 *  Use the next several functions to set the signals needed to
 *  load various registers
**/
function void loadPC(pcmux::pcmux_sel_t sel);
    load_pc = 1'b1;
    pcmux_sel = sel;
endfunction

function void loadRegfile(regfilemux::regfilemux_sel_t sel);
endfunction

function void loadMAR(marmux::marmux_sel_t sel);
endfunction

function void loadMDR();
endfunction

function void setALU(alumux::alumux1_sel_t sel1, alumux::alumux2_sel_t sel2, logic setop, alu_ops op);
    /* Student code here */


    if (setop)
        aluop = op; // else default value
endfunction

function automatic void setCMP(cmpmux::cmpmux_sel_t sel, branch_funct3_t op);
endfunction

/*****************************************************************************/

    /* Remember to deal with rst signal */
always_comb
begin : state_actions
    /* Default output assignments */
    set_defaults();
    /* Actions for each state */
    unique case(state)//?? some of these might take multiple clock cycles to complete

        f1: begin
            marmux_sel = marmux::pc_out;
            load_mar = 1'b1;
        end

        f2: begin
            mem_read = 1'b1;
            if(mem_resp)
                load_mdr = 1'b1;
            else 
                load_mdr = 1'b0;
        end

        f3: begin
            load_ir = 1'b1;
        end

        de: begin
            if((opcode == op_store) || (opcode == op_load)) begin //prime mar_o need it to determine how to shift rs2_out
                //load_data_out = 1'b1;
                marmux_sel = marmux::alu_out; //alu_out
                load_mar = 1'b1;
                alumux1_sel = alumux::rs1_out; //rs1
                alumux2_sel = alumux::s_imm; //s_imm
                $cast(alu_oppy, 3'b000); //add
                aluop = alu_oppy; 
            end
            else ;
        end

        imm: begin//need setup alu operands and control signals
            case(funct3)
                3'b000: begin   //addi
                    $cast(alu_oppy, 3'b000); //add
                    aluop = alu_oppy;
                    alumux1_sel = alumux::rs1_out; //rs1
                    alumux2_sel = alumux::i_imm; //i_imm
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::alu_out; //alu_out
                end

                3'b001: begin   //slli
                    $cast(alu_oppy, 3'b001); //sll
                    aluop = alu_oppy;
                    alumux1_sel = alumux::rs1_out; //rs1
                    alumux2_sel = alumux::i_imm; //i_imm
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::alu_out; //alu_out
                end

                3'b010: begin   //slti
                    cmpop = 3'b100; //blt
                    cmpmux_sel = cmpmux::i_imm; //i_imm
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::br_en; //zext br_en
                end

                3'b011: begin   //sltui
                    cmpop = 3'b110; //bltu
                    cmpmux_sel = cmpmux::i_imm; //i_imm
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::br_en; //zext br_en
                end
                
                3'b100: begin   //xori
                    $cast(alu_oppy, 3'b100); //xor
                    aluop = alu_oppy;
                    alumux1_sel = alumux::rs1_out; //rs1
                    alumux2_sel = alumux::i_imm; //i_imm
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::alu_out; //alu_out
                end

                3'b101: begin   //srli/srai based on bit 30
                    if(funct7[5]) begin
                        $cast(alu_oppy, 3'b010); //sra
                        aluop = alu_oppy;
                    end
                    else begin
                        $cast(alu_oppy, 3'b101); //srl
                        aluop = alu_oppy;
                    end
                    alumux1_sel = alumux::rs1_out; //rs1
                    alumux2_sel = alumux::i_imm; //i_imm
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::alu_out; //alu_out
                end

                3'b110: begin   //ori
                    $cast(alu_oppy, 3'b110); //or
                    aluop = alu_oppy;
                    alumux1_sel = alumux::rs1_out; //rs1
                    alumux2_sel = alumux::i_imm; //i_imm
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::alu_out; //alu_out
                end

                3'b111: begin    //andi
                    $cast(alu_oppy, 3'b111); //and
                    aluop = alu_oppy;
                    alumux1_sel = alumux::rs1_out; //rs1
                    alumux2_sel = alumux::i_imm; //i_imm
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::alu_out; //alu_out
                end

                default: ;
            endcase
            pcmux_sel = pcmux::pc_plus4; //pc_plus4
            load_pc = 1'b1;
        end

        lui: begin
            load_regfile = 1'b1;
            regfilemux_sel = regfilemux::u_imm; //u_imm
            pcmux_sel = pcmux::pc_plus4; //pc_plus4
            load_pc = 1'b1;
        end

        br: begin
            case (funct3)
                3'b000: begin   //beq
                    cmpop = 3'b000;
                    cmpmux_sel = cmpmux::rs2_out;
                end
                3'b001: begin   //bne
                    cmpop = 3'b001;
                    cmpmux_sel = cmpmux::rs2_out;
                end
                3'b100: begin   //blt
                    cmpop = 3'b100;
                    cmpmux_sel = cmpmux::rs2_out;
                end
                3'b101: begin   //bge
                    cmpop = 3'b101;
                    cmpmux_sel = cmpmux::rs2_out;
                end
                3'b110: begin   //bltu
                    cmpop = 3'b110;
                    cmpmux_sel = cmpmux::rs2_out;
                end
                3'b111: begin   //bgeu
                    cmpop = 3'b111;
                    cmpmux_sel = cmpmux::rs2_out;
                end
                default: begin  //beq default?
                    cmpop = 3'b000; 
                    cmpmux_sel = cmpmux::rs2_out;
                end
            endcase
            if(br_en) begin
                $cast(alu_oppy, 3'b000); //add
                aluop = alu_oppy;
                alumux1_sel = alumux::pc_out; //pc_out
                alumux2_sel = alumux::b_imm; //b_imm
                pcmux_sel = pcmux::alu_out; //alu_out
                load_pc = 1'b1;
            end
            else begin
                pcmux_sel = pcmux::pc_plus4; //pc_plus4
                load_pc = 1'b1;
            end
        end

        auipc: begin
            $cast(alu_oppy, 3'b000); //add
            aluop = alu_oppy;
            alumux1_sel = alumux::pc_out; //pc_out
            alumux2_sel = alumux::u_imm; //u_imm
            load_regfile = 1'b1;
            regfilemux_sel = regfilemux::alu_out; //alu_out
            pcmux_sel = pcmux::pc_plus4; //pc_plus4
            load_pc = 1'b1;
        end

        calc_addr: begin //a bit redundant given mar is changed in decode stage to prep for calculating the data_out value
            if(opcode == op_store) begin
                load_data_out = 1'b1;
                marmux_sel = marmux::alu_out; //alu_out
                load_mar = 1'b1;
                alumux1_sel = alumux::rs1_out; //rs1
                alumux2_sel = alumux::s_imm; //s_imm
                $cast(alu_oppy, 3'b000); //add
                aluop = alu_oppy;        
            end
            else begin
                marmux_sel = marmux::alu_out; //alu_out
                load_mar = 1'b1;
                alumux1_sel = alumux::rs1_out; //rs1
                alumux2_sel = alumux::i_imm; //i_imm
                $cast(alu_oppy, 3'b000);//add
                aluop = alu_oppy;
            end
        end

        ld1: begin
            mem_byte_enable = rmask;
            if(mem_resp) begin
                load_mdr = 1'b1;
                mem_read = 1'b1;
            end
            else begin
                mem_read = 1'b1;
            end
        end

        ld2: begin
            load_regfile = 1'b1;
            pcmux_sel = pcmux::pc_plus4; //pc_plus4
            load_pc = 1'b1;
            case (funct3)
                3'b000: begin   //lb
                    regfilemux_sel = regfilemux::lb; //lb 
                end
                3'b001: begin   //lh
                    regfilemux_sel = regfilemux::lh; //lh
                end
                3'b010: begin   //lw
                    regfilemux_sel = regfilemux::lw; //lw
                end
                3'b100: begin   //lbu
                    regfilemux_sel = regfilemux::lbu; //lbu
                end
                3'b101: begin   //lhu
                    regfilemux_sel = regfilemux::lhu; //lhu
                end
                default: ;
            endcase
        end

        st1: begin
            mem_byte_enable = wmask;
            if(mem_resp) begin
                load_mdr = 1'b1;
                mem_write = 1'b1;
            end
            else begin
                mem_write =1'b1;
            end
        end

        st2: begin
            load_pc = 1'b1;
            pcmux_sel = pcmux::pc_plus4; //pc_plus4
        end

        reg0: begin
            case(funct3)
                3'b000: begin   //add/sub
                    if(funct7[5]) begin
                        $cast(alu_oppy, 3'b011); //sub
                        aluop = alu_oppy;
                    end
                    else begin
                        $cast(alu_oppy, 3'b000); //add
                        aluop = alu_oppy;
                    end
                    alumux1_sel = alumux::rs1_out; //rs1
                    alumux2_sel = alumux::rs2_out; //rs2
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::alu_out; //alu_out
                end
                3'b001: begin   //sll
                    $cast(alu_oppy, 3'b001); //sll
                    aluop = alu_oppy;
                    alumux1_sel = alumux::rs1_out; //rs1
                    alumux2_sel = alumux::rs2_out; //rs2
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::alu_out; //alu_out
                end
                3'b010: begin   //slt
                    cmpop = 3'b100; //blt
                    cmpmux_sel = cmpmux::rs2_out; //rs2
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::br_en; //zext br_en
                end
                3'b011: begin   //sltu
                    cmpop = 3'b110; //bltu
                    cmpmux_sel = cmpmux::rs2_out; //rs2
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::br_en; //zext br_en
                end
                3'b100: begin   //xor
                    $cast(alu_oppy, 3'b100); //xor
                    aluop = alu_oppy;
                    alumux1_sel = alumux::rs1_out; //rs1
                    alumux2_sel = alumux::rs2_out; //rs2
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::alu_out; //alu_out
                end
                3'b101: begin   //srl/sra
                    if(funct7[5]) begin
                        $cast(alu_oppy, 3'b010); //sra
                        aluop = alu_oppy;
                    end
                    else begin
                        $cast(alu_oppy, 3'b101); //srl
                        aluop = alu_oppy;
                    end
                    alumux1_sel = alumux::rs1_out; //rs1
                    alumux2_sel = alumux::rs2_out; //rs2
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::alu_out; //alu_out
                end
                3'b110: begin   //or
                    $cast(alu_oppy, 3'b110); //add
                    aluop = alu_oppy;
                    alumux1_sel = alumux::rs1_out; //rs1
                    alumux2_sel = alumux::rs2_out; //rs2
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::alu_out; //alu_out
                end
                3'b111: begin   //and
                    $cast(alu_oppy, 3'b111); //add
                    aluop = alu_oppy;
                    alumux1_sel = alumux::rs1_out; //rs1
                    alumux2_sel = alumux::rs2_out; //rs2
                    load_regfile = 1'b1;
                    regfilemux_sel = regfilemux::alu_out; //alu_out
                end
            endcase
            pcmux_sel = pcmux::pc_plus4;
            load_pc = 1'b1;
        end

        jal: begin
            load_regfile = 1'b1;
            regfilemux_sel = regfilemux::pc_plus4;
            $cast(alu_oppy, 3'b000); //add
            aluop = alu_oppy;
            alumux1_sel = alumux::pc_out; //pc_out
            alumux2_sel = alumux::j_imm; //j_imm
            pcmux_sel = pcmux::alu_out; //alu_out
            load_pc = 1'b1;
        end

        jalr: begin
            load_regfile = 1'b1;
            regfilemux_sel = regfilemux::pc_plus4;
            $cast(alu_oppy, 3'b000); //add
            aluop = alu_oppy;
            alumux1_sel = alumux::rs1_out; //rs1
            alumux2_sel = alumux::i_imm; //i_imm
            pcmux_sel = pcmux::alu_mod2; //alu_mod2
            load_pc = 1'b1;
        end
        default: ;
    endcase
end

always_comb
begin : next_state_logic
    /* Next state information and conditions (if any)
     * for transitioning between states */
    unique case(state)
        f1: next_states = f2;

        f2: begin
            if(mem_resp)
                next_states = f3;
            else
                next_states = f2;
        end

        f3: next_states = de;

        de: begin
            case(opcode)
                op_lui: next_states = lui;
                op_imm: next_states = imm;
                op_br: next_states = br;
                op_auipc: next_states = auipc;
                op_load: next_states = calc_addr;
                op_store: next_states = calc_addr;
                op_reg: next_states = reg0;
                op_jal: next_states = jal;
                op_jalr: next_states = jalr;
                default: next_states = f1;
            endcase
        end

        imm: next_states = f1;

        lui: next_states = f1;

        br: begin
            next_states = f1;
        end

        auipc: next_states = f1;

        calc_addr: begin
            if(opcode == op_load)
                next_states = ld1;
            else
                next_states = st1; 
        end

        ld1: begin
            if(mem_resp)
                next_states = ld2;
            else
                next_states = ld1;
        end

        ld2: next_states = f1;

        st1: begin
            if(mem_resp)
                next_states = st2;
            else
                next_states = st1;
        end

        st2: next_states = f1;

        reg0: next_states = f1;

        jal: next_states = f1;

        jalr: next_states = f1;

        default: next_states = f1;
    endcase
end

always_ff @(posedge clk)
begin: next_state_assignment
    /* Assignment of next state on clock edge */
    if(rst)
        state <= f1;
    else
        state <= next_states;
end

endmodule : control
