package rv32i_cache_types;

typedef rv32i_word [7:0] rv32i_cacheline;

endpackage
